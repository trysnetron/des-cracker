------------------------------------------------
-------------------DES sim----------------------
------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.des_pkg.all;


entity des_sim is

end entity des_sim;


architecture sim of des_sim is

end architecture sim;
