
use work.des_pkg.all;


entity des_sim is

end entity des_sim;


architecture sim of des_sim is

end architecture sim;